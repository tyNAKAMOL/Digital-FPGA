// Verilog test fixture created from schematic E:\2D\Digital\finalAssignment\Final_Assignment_Digital_SmartHome\Counter_Up_0_3.sch - Wed Dec 15 11:33:49 2021

`timescale 1ns / 1ps

module Counter_Up_0_3_Counter_Up_0_3_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   Counter_Up_0_3 UUT (
		
   );
// Initialize Inputs
   initial begin
	CLK_IN = 0;
	end
endmodule
